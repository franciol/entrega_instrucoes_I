LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY UCONTROLE IS
    GENERIC (
        DATA_SIZE : NATURAL := 32
    );
    PORT (
        DATA : IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
        SAIDA_ULA : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		  SAIDA_PC, SAIDA_REG, SAIDA_MUXREG, SAIDA_MUXULA, SAIDA_MUXLOAD, SAIDA_MUXBEQ : OUT STD_LOGIC
    );
END ENTITY;

ARCHITECTURE arch OF UCONTROLE IS
BEGIN
    SAIDA_MUXBEQ <= "0" WHEN DATA(31 DOWNTO 26) = "000000" ELSE "1";  -- INSTRUCAO I RECEBE 1
	 SAIDA_MUXLOAD <= "0" WHEN DATA(31 DOWNTO 26) = "000000" ELSE "1";  -- INSTRUCAO I RECEBE 1
    SAIDA_MUXREG <= "0" WHEN DATA(31 DOWNTO 26) = "000000" ELSE "1";  -- INSTRUCAO I RECEBE 1
	 SAIDA_MUXULA <= "0" WHEN DATA(31 DOWNTO 26) = "000000" ELSE "1";  -- INSTRUCAO I RECEBE 1
    SAIDA_ULA <= "001" WHEN (DATA(31 DOWNTO 26) = "000000" AND DATA(5 DOWNTO 0) = "100000") ELSE
     ("010") WHEN (DATA(31 DOWNTO 26) = "000000" AND DATA(5 DOWNTO 0) = "100010") ELSE 
     ("000");
    

END arch;