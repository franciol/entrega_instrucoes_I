LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY UCONTROLE IS
    GENERIC (
        DATA_SIZE : NATURAL := 32
    );
    PORT (
        DATA : IN STD_LOGIC_VECTOR(DATA_SIZE-1 DOWNTO 0);
        SAIDA_PC, SAIDA_REG : OUT STD_LOGIC;
        SAIDA_ULA : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch OF UCONTROLE IS
BEGIN
    SAIDA_ULA <= DATA(5 DOWNTO 0) WHEN (DATA()) ELSE
END arch;